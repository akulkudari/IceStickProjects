module trafficcontroller(
    input clk_in, east_street, west_street
    
);

endmodule